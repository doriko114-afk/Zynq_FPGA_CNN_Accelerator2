`timescale 1ns / 1ps

module fc_layer #(
    parameter DATA_WIDTH = 20,
    parameter NUM_INPUTS = 676 // 13 * 13 * 4
)(
    input wire clk,
    input wire rst_n,
    input wire en,
    input wire valid_in,
    
    // �ǽð� ���� ����ġ �Է� (System Top���� 0 �Է� ��)
    input wire signed [31:0] adj_bias_0,
    input wire signed [31:0] adj_bias_1,
    input wire signed [31:0] adj_bias_2,

    // 4ä�� �Է� ���� ����
    input wire signed [DATA_WIDTH-1:0] data_in_0,
    input wire signed [DATA_WIDTH-1:0] data_in_1,
    input wire signed [DATA_WIDTH-1:0] data_in_2,
    input wire signed [DATA_WIDTH-1:0] data_in_3,
    
    output reg valid_out,
    output reg signed [31:0] score0, score1, score2
);

    // =========================================================================
    // [����ġ ������] Python Hardcore Mode ��� (Target: I, O, W)
    // =========================================================================

    // Class 0: O (Circle)
    localparam signed [31:0] BIAS_0_BASE = -20;
    localparam signed [7:0] W_0 [0:675] = '{
          -2,  -4,   0,  -2,   0,  -1,   0,   0,   2,   2,   3,   4,   6,
          -2,   0,   0,   0,   0,  -3,   0,   0,   2,   4,   5,   4,   5,
          -2,  -4,  -3,  -4,  -3,  -1,   2,   1,   2,   5,   3,   5,   5,
          -1,  -3,  -3,  -4,  -6,  -2,   0,   3,   4,   3,   1,   4,   7,
           1,  -1,  -2,  -1,  -3,  -2,   3,   3,   1,   3,   5,   4,   5,
           5,   3,   1,  -1,  -4,  -4,   0,   0,   0,   3,   4,   6,   8,
           8,   4,   5,   0,  -1,  -8, -10,  -3,  -1,  -2,   3,   8,  11,
          10,   4,   5,   1,   1,   0,  -6,  -3,  -2,  -4,  -2,   4,   5,
           7,   7,   1,   1,   0,  -1,  -2,  -3,  -4,  -6,  -4,  -2,   5,
           8,   3,   1,   1,   2,   1,  -2,  -6,  -4,  -6,  -4,  -2,  -1,
           4,   3,   1,   3,  -1,  -2,  -2,  -3,  -5,  -6,  -5,  -6,   0,
           0,   1,  -1,   0,   0,   0,  -3,  -4,  -8,  -4,  -5,  -6,  -6,
           0,   2,  -3,   0,  -4,  -5,  -5,  -7,  -6,  -3,  -3,  -4,  -5,
           0,   1,   1,   0,  -2,  -4,  -4,  -3,  -4,  -7,  -4,  -4,  -3,
           3,   4,   3,   1,   0,  -3,  -3,  -3,  -5,  -4,  -2,  -3,   0,
           1,   0,   0,   0,  -1,  -5,  -5,  -5,  -5,  -4,  -2,  -1,   3,
           3,   3,   1,   0,   0,  -1,  -3,  -6,  -4,  -4,  -2,   0,   3,
           3,   4,   3,   0,  -2,   0,  -3,  -4,  -4,  -2,   3,   0,   5,
           5,   4,   4,  -1,  -2,  -6,  -5,  -6,  -3,  -2,   1,   6,   6,
           5,   4,   1,   0,  -1,  -9, -12,  -5,  -5,   0,   6,   4,   7,
           6,   3,   0,   0,  -1,  -6, -12,   0,  -1,  -1,   4,   5,   7,
           2,   0,  -1,  -2,  -3,  -6,  -9,  -5,  -3,  -3,   0,   9,   9,
          -1,  -3,  -3,  -2,  -5,  -7,  -9,  -4,  -2,  -1,   0,   2,   7,
          -1,  -3,  -3,  -3,  -5,  -7,  -6,  -4,  -1,   0,   1,   2,   9,
          -5,  -3,  -3,  -4,  -4,  -6,  -6,  -5,  -6,  -2,   0,   0,  -2,
          -5,  -5,  -2,  -7,  -8,  -9,  -8,  -9,  -8,  -7,  -3,  -2,  -2,
           5,   0,   2,   0,   2,   5,   3,   6,   1,   1,   0,   6,   2,
           3,   3,   1,   4,   4,   3,   4,   6,   3,   4,   2,   0,   1,
           1,   1,   0,   2,   3,   7,   6,   6,   3,   4,   0,   0,   0,
           2,   2,   0,   2,   3,   5,   9,   9,   5,   2,   0,   0,   2,
           3,   0,   3,   2,   3,   2,   8,   7,   4,   5,   0,  -1,   0,
           6,   3,   7,   2,   3,   5,   4,   4,   4,   1,   2,   5,   1,
           6,   4,   1,   0,   0,   1,  -4,  -3,   1,   1,   2,   3,   3,
           6,   2,   0,   0,   1,   0,   2,   2,   1,   2,  -3,   0,   2,
           0,  -4,  -4,   0,   0,   1,   6,   2,   3,   3,  -1,   0,  -3,
          -4,  -1,  -1,  -1,   4,   5,   5,   4,   2,   3,   0,  -1,  -1,
          -3,   0,  -2,   0,   5,   5,   6,   3,   4,   2,   2,   0,  -2,
          -5,   0,  -1,   2,   6,   6,   6,   6,   5,   6,   2,   4,  -2,
          -6,   0,   1,   0,   3,   3,   4,   2,   1,   1,   2,   0,  -4,
          -4,  -3,   0,   1,   3,   2,   2,   0,   3,   4,   1,   2,  -6,
          -3,  -1,   0,  -1,  -1,   6,   4,   3,   4,   2,   1,   0,   0,
           0,   1,   1,   1,   1,   7,   6,   4,   1,   0,   0,   2,  -1,
           4,   2,   1,   1,   4,   2,   4,   3,   1,  -1,  -2,  -1,   0,
           0,   0,   3,   0,   3,   0,   2,   5,   1,   0,   2,   0,   3,
           6,   3,   2,   2,   2,   4,   5,   4,   3,   3,   3,   2,   2,
          10,   6,   6,   2,  -4,  -6,  -4,  -3,  -2,   0,   1,   2,   6,
          13,   5,   3,   0,  -3,  -9,  -9, -10,  -4,  -1,   3,   6,   5,
           8,   3,   0,  -2,  -2,  -2,   0,   0,  -3,   0,   1,   4,   6,
           7,   0,  -2,  -4,  -5,  -2,  -4,   0,   0,  -1,   1,   3,   5,
           1,  -2,  -3,  -4,  -2,  -2,  -2,  -1,   0,   0,   1,   0,   0,
          -5,  -3,  -3,   0,   0,   1,   3,   1,   2,   1,   0,   1,   3,
          -7,  -2,  -1,  -3,  -2,   0,   0,   1,  -2,   1,   0,   1,  -2
    };

    // Class 1: W (Square/Zigzag)
    localparam signed [31:0] BIAS_1_BASE = -32;
    localparam signed [7:0] W_1 [0:675] = '{
           0,  -1,  -2,   0,  -6,  -7,  -7,  -8, -11,  -7,  -6,  -2,  -6,
           0,  -1,   0,  -1,  -2,  -4,  -5,  -3,  -5,  -5,  -4,  -4,  -6,
           5,   1,   0,   0,   1,   0,  -4,  -4,  -3,  -3,  -4,  -2,   0,
           6,   5,   0,   0,  -3,  -3,  -9,  -7,  -2,  -5,  -3,  -8,   0,
           5,   7,   3,   0,   0,  -4, -11,  -7,  -5,  -3,  -3,   0,   0,
           7,   4,   4,   1,  -2,   0,  -2,   0,   2,  -1,  -4,   2,   0,
           5,   5,   6,   1,   3,   4,   6,   5,   3,   0,   1,   2,   2,
           8,   0,   2,   2,   0,   2,   4,   5,   4,   5,   4,   1,   3,
           5,   1,   2,   0,   0,   0,   3,   4,   2,   2,   3,   0,   6,
           6,   0,   0,   1,   2,   1,   1,   0,   4,   2,   0,   1,   4,
           3,   3,   4,   3,   0,  -1,   0,   0,   4,   2,   3,   2,   4,
           7,   0,  -1,   1,   0,  -2,  -2,   1,   1,   1,   0,   2,   5,
           6,   2,   4,   2,   4,   0,  -1,   1,   2,   3,   3,   1,   1,
          -2,   0,  -2,  -2,   0,  -3,  -4,   1,   1,   4,   3,   2,   2,
          -1,   0,   0,   0,   0,   0,   0,   4,   3,   1,   2,   7,   2,
           0,  -1,   0,   0,   1,  -2,   1,   1,   0,   2,   4,   4,   4,
           0,   1,   0,   2,   0,  -2,  -5,   0,   1,   0,   3,   3,   6,
           0,   1,   1,   0,  -1,  -1,  -6,  -1,   0,   0,   3,   3,   2,
          -1,   2,   2,   0,   0,  -1,   0,   1,   0,   0,   5,   4,   6,
           3,   1,   5,   0,   3,   4,   5,   0,  -1,   1,   3,   2,   6,
           2,   1,   2,   1,   4,   5,   4,   2,   1,   1,   4,   2,   7,
           1,   4,   3,   2,   0,   3,   3,   1,   0,  -2,   1,   3,   7,
           1,  -1,   2,   3,   1,   3,   3,   0,   1,   0,   1,   1,   8,
           1,   3,   1,   2,   0,   0,   1,   1,   1,  -2,   0,   3,   3,
           2,   3,   1,   3,   1,  -2,   0,   2,   1,   0,   2,   4,   0,
           3,   2,   2,   5,   0,   0,   1,   2,   2,   1,   5,   3,   4,
          -5,  -5,  -2,  -3,  -2,  -7,  -5,  -7,  -7,  -6,  -3,  -5,  -2,
           2,  -2,  -2,  -4,  -5,  -8,  -7,  -7,  -6,  -5,  -1,  -3,  -1,
           0,  -1,  -4,  -5,  -6,  -6,  -7,  -8,  -5,  -5,  -5,  -2,  -1,
           1,  -1,  -1,  -7,  -6, -10, -15,  -9,  -9,  -7,  -1,   2,   3,
           6,   0,  -1,  -6,  -1,  -4,  -7,  -4,  -3,  -2,  -2,   0,   1,
           7,   4,   0,  -2,   0,   0,   0,   0,   3,  -2,   0,   2,   8,
          10,   7,   6,   5,   4,   6,   4,   5,   5,   4,   4,   6,   7,
          10,   8,   3,   3,   1,   2,   0,   2,   1,   3,   4,   6,   6,
           5,   2,   2,   2,   2,  -1,   0,   1,   0,   1,   4,   2,   4,
           1,   1,   0,   0,   0,   0,  -2,  -4,  -3,  -1,   0,   1,   5,
           5,   1,   0,  -2,  -4,  -5,  -6,  -7,  -3,   0,  -3,   0,   2,
           2,   4,  -1,  -2,  -5,  -5,  -8,  -8,  -5,  -5,  -5,   0,   0,
           2,  -1,   0,   0,  -6,  -4,  -6,  -5,  -4,  -1,  -1,  -2,  -3,
          -2,  -3,  -5,  -7, -10, -11, -16, -12, -11, -10,  -8,  -4,   0,
          -2,  -2,  -1,  -4,  -4,  -5,  -6,  -7,  -5,  -5,  -2,   0,   0,
          -1,  -2,  -1,  -2,  -7,  -9,  -6,  -6,  -5,  -3,  -2,  -1,   1,
           0,   1,  -3,  -2,  -4,  -8,  -7, -10,  -5,  -3,  -1,   0,   3,
           2,  -2,  -1,  -2,  -7,  -8,  -8,  -9,  -7,  -2,  -3,   0,   6,
           3,   1,  -1,  -3,  -2,  -2,  -3,  -3,  -1,  -1,  -2,   3,   5,
           5,   2,   1,   3,   1,   5,   2,   7,   3,   2,   0,   5,  10,
           7,   7,   3,   3,   5,   6,   9,   9,   8,   5,   3,   6,   7,
           5,   5,   1,   2,   4,   5,   4,   6,   4,   2,   4,   5,   1,
           7,   3,   1,   0,   0,   4,   6,   4,   0,  -1,   0,   1,   3,
           7,   0,   0,   0,  -1,  -1,   0,  -1,  -1,   0,   1,   0,   3,
           5,   4,   2,   0,  -1,  -2,  -3,  -3,  -4,  -4,   2,   1,   1,
           5,   1,   3,  -5,  -3,  -4,  -5,  -5,  -2,  -2,   0,   2,   2
    };

    // Class 2: I (Triangle/Line)
    localparam signed [31:0] BIAS_2_BASE = 37;
    localparam signed [7:0] W_2 [0:675] = '{
           4,   2,   1,   3,  12,   7,   9,   9,   6,   0,  -1,   2,   1,
           0,   0,   2,   0,   1,   4,   5,   5,   2,  -4,   1,   0,  -3,
          -4,  -2,   0,   1,   4,   2,   7,   1,   1,  -3,   1,  -2,  -6,
          -6,  -4,   0,   4,   5,   6,   6,   1,   0,  -1,  -2,   2,  -6,
          -8,  -4,  -2,   1,   4,   7,   7,   3,   2,   1,  -2,  -3,  -7,
         -14, -10,  -7,   0,   3,   3,   0,   1,  -3,  -2,  -1,  -7, -10,
         -20, -17,  -8,  -2,   0,   1,   2,   2,  -3,   0,  -4, -13, -16,
         -22, -16, -16,  -4,  -1,   0,   3,   3,   0,   1,   0,  -7, -13,
         -16, -10,  -8,  -4,   1,   0,   2,  -1,   0,   1,   2,   0, -11,
         -17,  -4,  -3,  -3,   1,   0,   0,   1,   2,   2,   3,   4,  -3,
          -8,  -7,  -5,  -3,  -3,   1,   3,   3,   3,   2,   2,   2,  -3,
          -7,  -4,  -3,  -2,  -2,   1,   0,   4,   1,   2,   4,   1,  -1,
          -6,  -7,  -6,  -1,  -1,   6,   3,   7,   3,   0,   2,   0,   0,
           5,   0,   1,   0,   3,   6,   9,   3,   0,  -1,   0,  -1,   3,
          -4,  -1,   1,   0,   2,   5,   4,   5,   1,   2,   0,   0,   0,
           1,   0,  -2,   0,   0,   3,   7,   6,   1,   3,  -1,  -2,  -8,
          -4,  -4,  -1,  -1,   4,   4,   7,   6,   5,   0,  -3,  -3, -12,
          -3,  -6,  -3,  -2,   1,   2,   3,   5,   1,   1,  -6,  -6, -16,
          -7,  -8,  -6,  -2,   1,   0,   4,   3,   3,  -1,  -8,  -9, -18,
         -12, -16,  -6,   0,   0,   4,   6,   4,   0,  -2,  -9, -17, -25,
         -16, -11,  -3,  -1,   0,   7,   4,   2,   0,  -3,  -8, -16, -25,
          -8,   0,  -3,   1,   0,   4,   4,   1,   0,  -1,  -3, -11, -18,
          -5,   0,   0,   3,   5,   4,   3,   6,   3,   0,   0,  -8, -16,
          -2,   0,   0,   2,   5,   5,   6,   6,   2,   0,   0,  -5, -12,
           1,  -1,   0,   2,   6,   8,   6,   6,   2,   0,   0,  -2,  -2,
           0,   3,   3,   3,   7,   7,   8,   4,   4,   4,   0,  -1,   2,
           0,   2,   0,   0,   0,   2,   2,   2,   1,   1,   1,   0,   2,
          -4,   2,   2,   1,   3,   2,   0,   3,   0,   2,   0,   1,   1,
          -3,   2,   1,   0,   1,   3,   2,   1,   3,   2,   3,   1,  -2,
          -4,   1,  -1,   1,   2,   1,   3,   4,   1,   0,   2,   0,  -1,
          -7,  -3,   0,   0,   2,  -2,  -6,  -4,  -1,   1,   1,   0,  -6,
         -17, -10,  -9,  -2,   0,  -1,  -5,  -6,  -3,  -3,  -3, -11, -13,
         -24, -15, -10,  -4,  -5,  -4,  -2,  -1,  -2,  -5,  -8, -11, -16,
         -18,  -5,  -4,  -1,  -5,  -7,  -4,  -7,  -5,  -2,  -6,  -3, -12,
          -6,   0,   2,  -2,  -3,  -6,  -6,  -6,  -6,  -4,   0,  -1,  -5,
           0,   0,  -1,   0,  -1,  -3,  -5,   0,  -3,  -4,  -2,   0,  -4,
          -4,   0,   1,  -1,  -3,   0,   0,  -1,  -1,  -3,   1,   0,  -2,
           1,  -2,   0,   2,  -2,   0,   0,   0,   0,  -1,  -1,  -1,   1,
           2,   3,   3,  -1,   0,   5,   3,   2,   4,  -2,   2,   0,   3,
           8,   9,   5,   6,   5,   9,   7,  10,   9,   5,   2,   2,   3,
           4,   1,   0,   3,   2,   4,   4,   2,   4,   2,   0,   0,   0,
           0,   0,   0,   0,   3,   1,   0,   2,   0,   0,   1,   1,   1,
          -5,  -4,   1,   0,   0,   1,   1,   3,   3,   2,   3,   0,  -1,
          -4,   1,  -2,   1,   0,   5,   3,   6,   2,   1,   3,  -2,  -6,
         -14,  -8,  -4,  -2,   0,   0,  -2,  -2,   1,   0,   0,  -3,  -7,
         -18, -12,  -7,  -5,  -2,   0,  -2,   0,   0,  -2,  -5, -11, -18,
         -23, -17,  -7,  -1,   0,   1,   0,   5,   0,  -3,  -3, -13, -21,
         -18, -11,  -2,  -2,  -1,  -4,  -5,  -2,  -5,  -3,  -3,  -9, -13,
         -12,  -5,   0,   0,   2,   2,   0,  -1,   0,   0,   1,   0, -10,
          -6,   1,   0,   4,   2,   0,   0,   1,   0,   1,  -5,  -1,  -5,
           2,   0,   2,   0,  -1,   0,   0,   3,   1,   0,  -5,  -3,   0,
           0,   3,  -3,   4,   1,   5,   3,   4,   2,   2,  -2,  -3,  -4
    };

    // =========================================================================
    // Core Logic (Matrix Multiplication)
    // =========================================================================
    wire signed [31:0] FINAL_BIAS_0 = BIAS_0_BASE + adj_bias_0;
    wire signed [31:0] FINAL_BIAS_1 = BIAS_1_BASE + adj_bias_1;
    wire signed [31:0] FINAL_BIAS_2 = BIAS_2_BASE + adj_bias_2;

    reg signed [31:0] sum0, sum1, sum2;
    reg [9:0] counter; // 0 ~ 168 (169 pixels)
    reg processing;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            sum0 <= 0; sum1 <= 0; sum2 <= 0;
            counter <= 0; processing <= 0; valid_out <= 0;
        end else if (en && valid_in) begin
            if (!processing) begin
                // ù��° �ȼ� ���: �⺻ BIAS + ��ư ������(FINAL_BIAS) + 4ä�� ����
                // W Index mapping: Ch0(0~168), Ch1(169~337), Ch2(338~506), Ch3(507~675)
                sum0 <= FINAL_BIAS_0 + (data_in_0 * W_0[0]) + (data_in_1 * W_0[169]) + (data_in_2 * W_0[338]) + (data_in_3 * W_0[507]);
                sum1 <= FINAL_BIAS_1 + (data_in_0 * W_1[0]) + (data_in_1 * W_1[169]) + (data_in_2 * W_1[338]) + (data_in_3 * W_1[507]);
                sum2 <= FINAL_BIAS_2 + (data_in_0 * W_2[0]) + (data_in_1 * W_2[169]) + (data_in_2 * W_2[338]) + (data_in_3 * W_2[507]);
                counter <= 1; 
                processing <= 1;
                valid_out <= 0;
            end else begin
                // ���� ����
                sum0 <= sum0 + (data_in_0 * W_0[counter]) + (data_in_1 * W_0[counter+169]) + (data_in_2 * W_0[counter+338]) + (data_in_3 * W_0[counter+507]);
                sum1 <= sum1 + (data_in_0 * W_1[counter]) + (data_in_1 * W_1[counter+169]) + (data_in_2 * W_1[counter+338]) + (data_in_3 * W_1[counter+507]);
                sum2 <= sum2 + (data_in_0 * W_2[counter]) + (data_in_1 * W_2[counter+169]) + (data_in_2 * W_2[counter+338]) + (data_in_3 * W_2[counter+507]);
                
                if (counter == 168) begin // 169��° �ȼ�(�ε��� 168) ó�� �Ϸ�
                    processing <= 0;
                    valid_out <= 1;
                    score0 <= sum0; score1 <= sum1; score2 <= sum2;
                    counter <= 0;
                end else begin
                    counter <= counter + 1;
                end
            end
        end else valid_out <= 0;
    end
endmodule