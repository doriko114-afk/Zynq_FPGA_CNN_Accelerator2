------------------------------------------------------------------------------------
---- Engineer: Mike Field <hamster@snap.net.nz>
---- 
---- Description: Captures the pixels coming from the OV7670 camera and 
----              Stores them in block RAM
----
---- The length of href last controls how often pixels are captive - (2 downto 0) stores
---- one pixel every 4 cycles.
----
---- "line" is used to control how often data is captured. In this case every forth 
---- line
------------------------------------------------------------------------------------
--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

--entity ov7670_capture is
--    Port ( pclk  : in   STD_LOGIC;
--           rez_160x120 : IN std_logic;
--           rez_320x240 : IN std_logic;
--           sw    : in   STD_LOGIC_VECTOR(1 downto 0); -- [�߰�] ����ġ �Է�
--           vsync : in   STD_LOGIC;
--           href  : in   STD_LOGIC;
--           d     : in   STD_LOGIC_VECTOR (7 downto 0);
--           addr  : out  STD_LOGIC_VECTOR (18 downto 0);
--           dout  : out  STD_LOGIC_VECTOR (11 downto 0);
--           we    : out  STD_LOGIC);
--end ov7670_capture;

--architecture Behavioral of ov7670_capture is
--   signal d_latch      : std_logic_vector(15 downto 0) := (others => '0');
--   signal address      : STD_LOGIC_VECTOR(18 downto 0) := (others => '0');
--   signal line         : std_logic_vector(1 downto 0)  := (others => '0');
--   signal href_last    : std_logic_vector(6 downto 0)  := (others => '0');
--   signal we_reg       : std_logic := '0';
--   signal href_hold    : std_logic := '0';
--   signal latched_vsync : STD_LOGIC := '0';
--   signal latched_href  : STD_LOGIC := '0';
--   signal latched_d     : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
--begin

--	addr <= address;
--	we <= we_reg;
----	dout <= d_latch(15 downto 12) & d_latch(10 downto 7) & d_latch(4 downto 1); 
   
--	capture_process: process(pclk)
--	begin
--		if rising_edge(pclk) then
--			if we_reg = '1' then
--				address <= std_logic_vector(unsigned(address)+1);
--			end if;

--			-- This is a bit tricky href starts a pixel transfer that takes 3 cycles
--			--        Input   | state after clock tick   
--			--         href   | wr_hold    d_latch           dout                we address  address_next
--			-- cycle -1  x    |    xx      xxxxxxxxxxxxxxxx  xxxxxxxxxxxx  x   xxxx     xxxx
--			-- cycle 0   1    |    x1      xxxxxxxxRRRRRGGG  xxxxxxxxxxxx  x   xxxx     addr
--			-- cycle 1   0    |    10      RRRRRGGGGGGBBBBB  xxxxxxxxxxxx  x   addr     addr
--			-- cycle 2   x    |    0x      GGGBBBBBxxxxxxxx  RRRRGGGGBBBB  1   addr     addr+1

--			-- detect the rising edge on href - the start of the scan line
--			if href_hold = '0' and latched_href = '1' then
--				case line is
--					when "00"   => line <= "01";
--					when "01"   => line <= "10";
--					when "10"   => line <= "11";
--					when others => line <= "00";
--				end case;
--			end if;
--			href_hold <= latched_href;
         
--			-- capturing the data from the camera, 12-bit RGB
--			if latched_href = '1' then
--				d_latch <= d_latch( 7 downto 0) & latched_d;
--			end if;
--			we_reg  <= '0';

--			-- Is a new screen about to start (i.e. we have to restart capturing
--			if latched_vsync = '1' then 
--				address      <= (others => '0');
--				href_last    <= (others => '0');
--				line         <= (others => '0');
--			else
--                -- (1) ���� Ÿ�̹� ����: href_last�� 0�� ��Ʈ�� 1�� �� (2Ŭ������ 1����)
--                if href_last(0) = '1' then 
                    
--                    we_reg <= '1';                -- �޸𸮿� ���� ���
--                    href_last <= (others => '0'); -- Ÿ�̹� ����

--                    -- (2) ������ ���� (YUV ����� ����)
--                    -- YUV ��忡�� d�� Y/U/V�� ���� ���ɴϴ�.
--                    -- ���� ��ü�� V���� �ſ� �����Ƿ�(���� 140~150 �̻�), 
--                    -- ������ ������(d)�� �ռ� ������(latched_d) �� �ϳ��� ũ�� ������� ǥ���մϴ�.
                    
--                    case sw is
--                        when "00" => -- [������ ���] V���� ������ �˻�
--                            if unsigned(d) > 160 then
--                                dout <= x"FFF"; -- ��� (Ž����)
--                            else
--                                dout <= x"000"; -- ������
--                            end if;
                            
--                        when "01" => -- [�Ķ��� ���] U���� ������ �˻�
--                             -- �Ķ��� ��ü�� U���� ���� ���ɴϴ�.
--                             -- (����: YUV raw stream������ U�� V�� ���� ���� �˻��ϹǷ� 
--                             -- ������ ��ü�� ������ �� ������, �Ķ� ��ü�� ��� �� �νĵ˴ϴ�)
--                            if unsigned(d) > 150 then 
--                                dout <= x"FFF"; 
--                            else
--                                dout <= x"000"; 
--                            end if;
                            
--                        when "10" => -- [�ʷϻ� ���] V/U ���� ������ �˻�
--                            -- �ʷϻ��� U, V ������ ��� �����ϴ�.
--                            -- ��, ������(��ο� ��)�� ���� �����Ƿ�, �ʹ� ��ο� �� �����ؾ� �մϴ�.
--                            -- ����: ����(d)�� ����(90����) AND ���� ������(���, latched_d)�� ������ ��ƾ� ��(60�̻�)
--                            if (unsigned(d) < 90) and (unsigned(latched_d) > 60) then
--                                dout <= x"FFF";
--                            else
--                                dout <= x"000";
--                            end if;
                            
--                        when others => -- [��Ÿ: 11] �׳� ����ó�� �����Ű�ų� ������
--                             dout <= x"000";
--                    end case;

--                else
--                    -- Ÿ�̹��� �� ���� ���� �����͸� ����Ʈ�ϸ� ���
--                    we_reg <= '0';
--                    href_last <= href_last(href_last'high-1 downto 0) & latched_href;
--                end if;
--            end if;
                
--		end if;
	  
--		if falling_edge(pclk) then
--			latched_d     <= d;
--			latched_href  <= href;
--			latched_vsync <= vsync;
--		end if;	  
--	end process;
--end Behavioral;

--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

--entity ov7670_capture is
--    Port ( pclk  : in   STD_LOGIC;
--           rez_160x120 : IN std_logic; -- ��Ʈ�� �����ϵ� ���ο��� ����
--           rez_320x240 : IN std_logic; -- ��Ʈ�� �����ϵ� ���ο��� ����
--           sw    : in   STD_LOGIC_VECTOR(1 downto 0);
--           btn_up   : in STD_LOGIC;
--           btn_down : in STD_LOGIC;
--           vsync : in   STD_LOGIC;
--           href  : in   STD_LOGIC;
--           d     : in   STD_LOGIC_VECTOR (7 downto 0);
--           addr  : out  STD_LOGIC_VECTOR (18 downto 0);
--           dout  : out  STD_LOGIC_VECTOR (11 downto 0);
--           we    : out  STD_LOGIC;
--           x_center : out STD_LOGIC_VECTOR(9 downto 0);
--           y_center : out STD_LOGIC_VECTOR(9 downto 0)
--           );
--end ov7670_capture;

--architecture Behavioral of ov7670_capture is
--   signal d_latch      : std_logic_vector(15 downto 0) := (others => '0');
--   signal address      : STD_LOGIC_VECTOR(18 downto 0) := (others => '0');
--   signal href_last    : std_logic_vector(6 downto 0)  := (others => '0');
--   signal we_reg       : std_logic := '0';
--   signal latched_vsync : STD_LOGIC := '0';
--   signal latched_href  : STD_LOGIC := '0';
--   signal latched_d     : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');

--   -- �����߽� ��� ����
--   signal sum_x : unsigned(31 downto 0) := (others => '0');
--   signal sum_y : unsigned(31 downto 0) := (others => '0');
--   signal pixel_cnt : unsigned(19 downto 0) := (others => '0');
--   signal x_curr : unsigned(9 downto 0) := (others => '0');
--   signal y_curr : unsigned(9 downto 0) := (others => '0');
--   signal x_result : std_logic_vector(9 downto 0) := (others => '0');
--   signal y_result : std_logic_vector(9 downto 0) := (others => '0');

--   -- �Ӱ谪 (�ʱⰪ 50)
--   signal threshold_val : unsigned(19 downto 0) := to_unsigned(50, 20);

--begin
--   addr <= address;
--   we <= we_reg;
--   x_center <= x_result;
--   y_center <= y_result;
   
--   capture_process: process(pclk)
--   begin
--      if rising_edge(pclk) then
--         -- [����] �ػ� ������� ���� ��ȣ ������ ������ �ּ� ����
--         if we_reg = '1' then
--            address <= std_logic_vector(unsigned(address)+1);
--         end if;

--         -- href_last�� Ÿ�̹� ���߱�� ����Ʈ ��������
--         -- OV7670�� �⺻������ YUV/RGB �����͸� 2Ŭ���� 1�ȼ�(2����Ʈ) ����
         
--         -- ������ ��ġ (���� ����Ʈ + ���� ����Ʈ ���տ�)
--         if latched_href = '1' then
--            d_latch <= d_latch( 7 downto 0) & latched_d;
--         end if;
--         we_reg  <= '0';

--         -- VSYNC: ������ ����
--         if latched_vsync = '1' then 
--            address      <= (others => '0');
--            href_last    <= (others => '0');
--            x_curr <= (others => '0');
--            y_curr <= (others => '0');

--            -- ��ư���� �Ӱ谪 ����
--            if btn_up = '1' then
--                if threshold_val < 50000 then threshold_val <= threshold_val + 50; end if;
--            elsif btn_down = '1' then
--                if threshold_val > 50 then threshold_val <= threshold_val - 50; end if;
--            end if;

--            -- �����߽� ��� ��� ������Ʈ
--            if pixel_cnt > threshold_val then
--               x_result <= std_logic_vector(resize(sum_x / pixel_cnt, 10));
--               y_result <= std_logic_vector(resize(sum_y / pixel_cnt, 10));
--            end if;

--            sum_x <= (others => '0');
--            sum_y <= (others => '0');
--            pixel_cnt <= (others => '0');
         
--         else
--            -- VSYNC �ƴ� �� ������ ó��
            
--            -- [����] HREF�� Rising Edge�� �� (�� ���� ����) -> Y��ǥ ����
--            -- latched_href�� 0->1�� ���ϴ� ������ �����ϴ� ������ �ʿ�������
--            -- ���⼭�� ������ href_last ��Ʈ�� �̿��ϰų� href ��ȣ ��ü�� ���ϴ�.
--            -- ���� ������ �ܼ�ȭ: href�� 0�̾��ٰ� 1�� �Ǵ� ������ y_curr ���� �ʿ�
            
--            -- (����ȭ�� Y ���� ����)
--            -- href�� Low���ٰ� High�� �ö���� ���� üũ�� ���� �����ϹǷ�,
--            -- ���⼭�� x_curr�� 639(�� �� ��)�� �����ϸ� y_curr�� �ø��� ��� ���
            
--            if href_last(0) = '1' then 
--               we_reg <= '1';
--               href_last <= (others => '0');
               
--               x_curr <= x_curr + 1;
--               if x_curr = 639 then -- 640��° �ȼ��̸�
--                  x_curr <= (others => '0');
--                  y_curr <= y_curr + 1;
--               end if;

--               -- ���� ��� �� ���͸�
--               dout <= x"000"; 
               
--               case sw is
--                  when "00" => -- ����
--                     if unsigned(d) > 160 then
--                        dout <= x"FFF";
--                        sum_x <= sum_x + x_curr;
--                        sum_y <= sum_y + y_curr;
--                        pixel_cnt <= pixel_cnt + 1;
--                     end if;
--                  when "01" => -- �Ķ�
--                     if unsigned(d) > 160 then
--                        dout <= x"FFF";
--                        sum_x <= sum_x + x_curr;
--                        sum_y <= sum_y + y_curr;
--                        pixel_cnt <= pixel_cnt + 1;
--                     end if;
--                  when "10" => -- �ʷ�
--                     if (unsigned(d) < 80) and (unsigned(latched_d) > 60) then
--                        dout <= x"FFF";
--                        sum_x <= sum_x + x_curr;
--                        sum_y <= sum_y + y_curr;
--                        pixel_cnt <= pixel_cnt + 1;
--                     end if;
--                  when others => 
--                     -- �Ϲ� ���� (RGB444)
--                     dout <= d_latch(15 downto 12) & d_latch(10 downto 7) & d_latch(4 downto 1);
--               end case;

--            else
--               we_reg <= '0';
--               href_last <= href_last(href_last'high-1 downto 0) & latched_href;
--            end if;
--         end if;
--      end if;
      
--      if falling_edge(pclk) then
--         latched_d     <= d;
--         latched_href  <= href;
--         latched_vsync <= vsync;
--      end if;     
--   end process;
--end Behavioral;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ov7670_capture is
    Port ( pclk  : in   STD_LOGIC;
           rez_160x120 : IN std_logic;
           rez_320x240 : IN std_logic;
           sw    : in   STD_LOGIC_VECTOR(1 downto 0);
           btn_up   : in STD_LOGIC;
           btn_down : in STD_LOGIC;
           vsync : in   STD_LOGIC;
           href  : in   STD_LOGIC;
           d     : in   STD_LOGIC_VECTOR (7 downto 0);
           addr  : out  STD_LOGIC_VECTOR (18 downto 0);
           dout  : out  STD_LOGIC_VECTOR (11 downto 0);
           we    : out  STD_LOGIC;
           x_center : out STD_LOGIC_VECTOR(9 downto 0);
           y_center : out STD_LOGIC_VECTOR(9 downto 0)
           );
end ov7670_capture;

architecture Behavioral of ov7670_capture is
   signal d_latch      : std_logic_vector(15 downto 0) := (others => '0');
   signal address      : STD_LOGIC_VECTOR(18 downto 0) := (others => '0');
   signal href_last    : std_logic_vector(6 downto 0)  := (others => '0');
   signal we_reg       : std_logic := '0';
   signal latched_vsync : STD_LOGIC := '0';
   signal latched_href  : STD_LOGIC := '0';
   signal latched_d     : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
   
   -- �����߽� ��� ����
   signal sum_x : unsigned(31 downto 0) := (others => '0');
   signal sum_y : unsigned(31 downto 0) := (others => '0');
   signal pixel_cnt : unsigned(19 downto 0) := (others => '0');
   signal x_curr : unsigned(9 downto 0) := (others => '0');
   signal y_curr : unsigned(9 downto 0) := (others => '0');
   signal x_result : std_logic_vector(9 downto 0) := (others => '0');
   signal y_result : std_logic_vector(9 downto 0) := (others => '0');
   
   -- �Ӱ谪 (�ʱⰪ 50)
   signal threshold_val : unsigned(19 downto 0) := to_unsigned(50, 20);

begin
   addr <= address;
   we <= we_reg;
   x_center <= x_result;
   y_center <= y_result;
   
   capture_process: process(pclk)
   begin
      if rising_edge(pclk) then
         -- �ּ� ����
         if we_reg = '1' then
            address <= std_logic_vector(unsigned(address)+1);
         end if;

         -- ������ ��ġ
         if latched_href = '1' then
            d_latch <= d_latch( 7 downto 0) & latched_d;
         end if;
         we_reg  <= '0';

         -- VSYNC: ������ ����
         if latched_vsync = '1' then 
            address      <= (others => '0');
            href_last    <= (others => '0');
            x_curr <= (others => '0');
            y_curr <= (others => '0');
            
            -- ��ư���� �Ӱ谪 ����
            if btn_up = '1' then
                if threshold_val < 50000 then threshold_val <= threshold_val + 50; end if;
            elsif btn_down = '1' then
                if threshold_val > 50 then threshold_val <= threshold_val - 50; end if;
            end if;

            -- �����߽� ��� ������Ʈ
            if pixel_cnt > threshold_val then
               x_result <= std_logic_vector(resize(sum_x / pixel_cnt, 10));
               y_result <= std_logic_vector(resize(sum_y / pixel_cnt, 10));
            end if;

            sum_x <= (others => '0');
            sum_y <= (others => '0');
            pixel_cnt <= (others => '0');
         
         else
            -- VSYNC �ƴ� ��
            if href_last(0) = '1' then 
               we_reg <= '1';
               href_last <= (others => '0');
               
               -- ��ǥ ����
               x_curr <= x_curr + 1;
               if x_curr = 639 then 
                  x_curr <= (others => '0');
                  y_curr <= y_curr + 1;
               end if;

               -- [���� �Ϸ�] �ϴ� ������ ���͸� (Y��ǥ�� 478���� ���� ���� �ν�)
               dout <= x"000"; -- �⺻ ������
               
               if (y_curr < 478) then -- **478�� ������** (477 ���α��� ��ȿ)
                   case sw is
                      when "00" => -- ���� ����
                         if unsigned(d) > 160 then
                            dout <= x"FFF";
                            sum_x <= sum_x + x_curr;
                            sum_y <= sum_y + y_curr;
                            pixel_cnt <= pixel_cnt + 1;
                         end if;
                      when "01" => -- �Ķ� ����
                         if unsigned(d) > 160 then
                            dout <= x"FFF";
                            sum_x <= sum_x + x_curr;
                            sum_y <= sum_y + y_curr;
                            pixel_cnt <= pixel_cnt + 1;
                         end if;
                      when "10" => -- �ʷ� ����
                         if (unsigned(d) < 80) and (unsigned(latched_d) > 60) then
                            dout <= x"FFF";
                            sum_x <= sum_x + x_curr;
                            sum_y <= sum_y + y_curr;
                            pixel_cnt <= pixel_cnt + 1;
                         end if;
                      when others => 
                         -- �Ϲ� ����
                         dout <= d_latch(15 downto 12) & d_latch(10 downto 7) & d_latch(4 downto 1);
                   end case;
               end if; 
               
            else
               we_reg <= '0';
               href_last <= href_last(href_last'high-1 downto 0) & latched_href;
            end if;
         end if;
      end if;
      
      if falling_edge(pclk) then
         latched_d     <= d;
         latched_href  <= href;
         latched_vsync <= vsync;
      end if;     
   end process;
end Behavioral;