`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/07/06 21:38:58
// Design Name: 
// Module Name: ov7670_registers_2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ov7670_registers_2(
    input clk,  //50MHz clk �ޱ�
    input resend,  //debouce���� ���ΰ�ħ�ϴ� ���� �ޱ�
    input advance,  //���ΰ�ħ�� ������� �ϴ� ���� ����
    output [15:0] command,  // OV7670�� ���� �������� �� �� ������
    output finished  //������ �Ϸ�Ǿ����� ��Ÿ���� ��ȣ
);

    //���� ��ȣ
    reg [15:0] sreg;  //�������� �ּҸ� ��Ÿ���� ����
    reg finished_temp;  //������ �Ϸ�Ǿ����� ��Ÿ���� ��ȣ
    reg [7:0] address = {8{1'b0}};  //�ּ��� ũ��� �˳��� 8��Ʈ
    
    //��¿� �� �Ҵ�
    assign command = sreg;  // OV7670�� ���� �������� �� �� �����͸� Conroller���� ����ϴ� command ������ �ű�
    assign finished = finished_temp;  //������ �Ϸ�Ǿ����� ��Ÿ���� ��ȣ�� Conroller���� ����ϴ� finished ������ �ű�
    
    //�������Ϳ� ���� FFFF �� ���
    //������ �Ϸ�Ǿ����� ��Ÿ���� ��ȣ�� ǥ�õ˴ϴ�.(finished_temp)
    always @ (sreg) begin
        if(sreg == 16'hFFFF) begin
            finished_temp <= 1;
        end
        else begin
            finished_temp <= 0;  //������ �Ϸ���� �ʾҴ�.
        end
    end
    
    //lookuptable���� ������ ���(�������Ϳ���)
    always @ (posedge clk) begin
        if(resend == 1) begin           //���ΰ�ħ ��ȣ
            address <= {8{1'b0}};       //�ʱ�ȭ
        end
        else if(advance == 1) begin     //�ƴ϶�� ���� ������ ���
            address <= address+1;       //�ּҰ��� 1�� �����ָ鼭 ���ϴ� �������� ���� ã��
        end
           
        case (address)  //�ּ��� ���� ���� ���ϴ� �������Ϳ� ���� ���� ������ ����(�� �������� i2c����� ���)
                0:  sreg <= 16'h12_80; //reset
                1:  sreg <= 16'hFF_F0; //delay
                2:  sreg <= 16'h12_00; // COM7,     set RGB color output
                3:  sreg <= 16'h11_80; // CLKRC     internal PLL matches input clock
                4:  sreg <= 16'h0C_00; // COM3,     default settings
                5:  sreg <= 16'h3E_00; // COM14,    no scaling, normal pclock
                6:  sreg <= 16'h04_00; // COM1,     disable CCIR656
                7:  sreg <= 16'h40_d0; //COM15,     RGB565, full output range
                8:  sreg <= 16'h3a_04; //TSLB       set correct output data sequence (magic)
                9:  sreg <= 16'h14_18; //COM9       MAX AGC value x4
                10: sreg <= 16'h4F_B3; //MTX1       all of these are magical matrix coefficients
                11: sreg <= 16'h50_B3; //MTX2
                12: sreg <= 16'h51_00; //MTX3
                13: sreg <= 16'h52_3d; //MTX4
                14: sreg <= 16'h53_A7; //MTX5
                15: sreg <= 16'h54_E4; //MTX6
                16: sreg <= 16'h58_9E; //MTXS
                17: sreg <= 16'h3D_C0; //COM13      sets gamma enable, does not preserve reserved bits, may be wrong?
                18: sreg <= 16'h17_14; //HSTART     start high 8 bits
                19: sreg <= 16'h18_02; //HSTOP      stop high 8 bits //these kill the odd colored line
                20: sreg <= 16'h32_80; //HREF       edge offset
                21: sreg <= 16'h19_03; //VSTART     start high 8 bits
                22: sreg <= 16'h1A_7B; //VSTOP      stop high 8 bits
                23: sreg <= 16'h03_0A; //VREF       vsync edge offset
                24: sreg <= 16'h0F_41; //COM6       reset timings
                25: sreg <= 16'h1E_00; //MVFP       disable mirror / flip //might have magic value of 03
                26: sreg <= 16'h33_0B; //CHLF       //magic value from the internet
                27: sreg <= 16'h3C_78; //COM12      no HREF when VSYNC low
                //28: sreg <= 16'h69_00; //GFIX       fix gain control
                28: sreg <= 16'h69_0a; //GFIX  
                29: sreg <= 16'h74_00; //REG74      Digital gain control
                30: sreg <= 16'hB0_84; //RSVD       magic value from the internet *required* for good color
                31: sreg <= 16'hB1_0c; //ABLC1
                32: sreg <= 16'hB2_0e; //RSVD       more magic internet values
                33: sreg <= 16'hB3_80; //THL_ST
                //begin mystery scaling numbers
                34: sreg <= 16'h70_3a;
                35: sreg <= 16'h71_35;
                36: sreg <= 16'h72_11;
                37: sreg <= 16'h73_f0;
                38: sreg <= 16'ha2_02;
                //gamma curve values
                39: sreg <= 16'h7a_20;
                40: sreg <= 16'h7b_10;
                41: sreg <= 16'h7c_1e;
                42: sreg <= 16'h7d_35;
                43: sreg <= 16'h7e_5a;
                44: sreg <= 16'h7f_69;
                45: sreg <= 16'h80_76;
                46: sreg <= 16'h81_80;
                47: sreg <= 16'h82_88;
                48: sreg <= 16'h83_8f;
                49: sreg <= 16'h84_96;
                50: sreg <= 16'h85_a3;
                51: sreg <= 16'h86_af;
                52: sreg <= 16'h87_c4;
                53: sreg <= 16'h88_d7;
                54: sreg <= 16'h89_e8;
                //AGC and AEC
                55: sreg <= 16'h13_e0; //COM8, disable AGC / AEC
                56: sreg <= 16'h00_00; //set gain reg to 0 for AGC
                57: sreg <= 16'h10_00; //set ARCJ reg to 0
                58: sreg <= 16'h0d_40; //magic reserved bit for COM4
                59: sreg <= 16'h14_18; //COM9, 4x gain + magic bit
                60: sreg <= 16'ha5_05; // BD50MAX
                61: sreg <= 16'hab_07; //DB60MAX
                62: sreg <= 16'h24_95; //AGC upper limit
                63: sreg <= 16'h25_33; //AGC lower limit
                64: sreg <= 16'h26_e3; //AGC/AEC fast mode op region
                65: sreg <= 16'h9f_78; //HAECC1
                66: sreg <= 16'ha0_68; //HAECC2
                67: sreg <= 16'ha1_03; //magic
                68: sreg <= 16'ha6_d8; //HAECC3
                69: sreg <= 16'ha7_d8; //HAECC4
                70: sreg <= 16'ha8_f0; //HAECC5
                71: sreg <= 16'ha9_90; //HAECC6
                72: sreg <= 16'haa_94; //HAECC7
                73: sreg <= 16'h13_e5; //COM8, enable AGC / AEC
                default : sreg <= 16'hFFFF;  //sreg���� ffff�̸� ������ �Ϸ� �Ǿ���.
        endcase
    end
endmodule

module ov7670_registers_setting_tb;

    reg clk=0;
    reg resend;
    reg advance=0;
    wire [15:0] command;
    wire finished;
    
    ov7670_registers_2 uut(clk, resend, advance, command, finished);
    
    always #10 clk=~clk; 
    initial begin
        #100 resend=1;
        #100 resend=0;
    end
    
    always #300 advance = ~advance;
    
endmodule