`timescale 1ns / 1ps
`default_nettype none

module cnn_top #(
    parameter IMG_WIDTH  = 28,  // �ùķ��̼�/�׽�Ʈ��
    parameter IMG_HEIGHT = 28,
    parameter DATA_WIDTH = 8,
    parameter FC_INPUTS  = 169
)(
    input wire clk,           // �ý��� Ŭ�� (��: 125MHz or 100MHz)
    input wire clk_pix,       // �ȼ� Ŭ�� (25MHz, Clock Wizard���� �����Ǿ� ����)
    input wire clk_tmds,      // HDMI ��� Ŭ�� (250MHz, Clock Wizard���� �����Ǿ� ����)
    input wire rst_n,
    
    // [�ٽ�] ����ġ �Է� (System Top���� ��������� ��)
    // sw[0]: ���̵���� �ڽ� ON/OFF
    // sw[1]: ��� ���� (Freeze)
    // sw[2]: CNN ���� ���� & �ؽ�Ʈ ��� ON
    input wire [2:0] sw,

    // ī�޶�/���� �Է�
    input wire cam_href,      // HSYNC ����
    input wire cam_vsync,     // VSYNC ����
    input wire [7:0] cam_data, // ���� ������ (Grayscale ����)

    // CNN�� ����ġ �Է� (���� ��⿡�� ����� �����ϰų� �������ͷ� ����)
    input wire signed [DATA_WIDTH-1:0] k00, k01, k02,
    input wire signed [DATA_WIDTH-1:0] k10, k11, k12,
    input wire signed [DATA_WIDTH-1:0] k20, k21, k22,
    input wire signed [DATA_WIDTH-1:0] bias,

    // HDMI ��� ��Ʈ
    output wire [2:0] tmds_data_p, tmds_data_n,
    output wire tmds_clk_p, tmds_clk_n,
    
    // ������ LED (���û���)
    output wire [2:0] led_check
);

    // =============================================================
    // 1. ���� ��ȣ ����
    // =============================================================
    wire conv_valid;
    wire signed [19:0] conv_data;
    
    wire class_valid;
    wire signed [31:0] score_c, score_t, score_s;
    
    // ��� ó����
    reg [1:0] current_winner;   // �ǽð� 1��
    reg [1:0] final_result;     // ���� ǥ�ÿ� (Freeze �����)
    reg [2:0] osd_msg_code;     // RGB ���� ���� �ڵ�

    // ���� ������ ó�� (8bit -> 12bit Ȯ��)
    wire [11:0] osd_din;
    assign osd_din = {cam_data[7:4], cam_data[7:4], cam_data[7:4]}; // ����� RGB��

    // =============================================================
    // 2. CNN ���� ��� (Conv -> FC)
    // =============================================================
    
    // (1) Conv Layer
    conv_layer_top #(
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        .DATA_WIDTH(DATA_WIDTH)
    ) u_conv_layer (
        .clk(clk),
        .rst_n(rst_n),
        .valid_in(cam_href),   // ���� ���� �� valid��� ���� (���� Ÿ�̹� �°� ���� �ʿ�)
        .data_in(cam_data),
        
        .k00(k00), .k01(k01), .k02(k02),
        .k10(k10), .k11(k11), .k12(k12),
        .k20(k20), .k21(k21), .k22(k22),
        .bias(bias),
        
        .valid_out(conv_valid),
        .layer_out(conv_data)
    );

    // (2) FC Layer (������ ���� ���)
    fc_layer #(
        .DATA_WIDTH(20),
        .NUM_INPUTS(FC_INPUTS)
    ) u_fc_layer (
        .clk(clk),
        .rst_n(rst_n),
        .en(sw[2]),            // SW2�� ������ ���� ����
        .valid_in(conv_valid),
        .data_in(conv_data),
        
        .valid_out(class_valid),
        .score0(score_c),
        .score1(score_t),
        .score2(score_s)
    );

    // =============================================================
    // 3. ��� �Ǵ� �� ����ġ ���� ���� (SW1 Freeze)
    // =============================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            final_result <= 0;
            current_winner <= 0;
            osd_msg_code <= 0;
        end else begin
            // A. ���� ������ ���� ���� ã��
            if (score_c >= score_t && score_c >= score_s) current_winner <= 2'd0; // ��
            else if (score_t >= score_c && score_t >= score_s) current_winner <= 2'd1; // �ﰢ��
            else current_winner <= 2'd2; // �簢��

            // B. SW1 (Freeze) ����
            if (sw[1] == 1'b0) begin
                // ����ġ ���� -> �ǽð� ��� �ݿ�
                final_result <= current_winner;
            end 
            // ����ġ ����(1) -> else�� �� �����ν� ���� �� ���� (Latch/Freeze)

            // C. RGB ���� �޽��� �ڵ�� ��ȯ
            case (final_result)
                2'd0: osd_msg_code <= 3'b001; // CIR
                2'd1: osd_msg_code <= 3'b010; // TRI
                2'd2: osd_msg_code <= 3'b011; // REC
                default: osd_msg_code <= 3'b000;
            endcase
        end
    end

    // LED�� ���� ����� (���� ���� ��������)
    assign led_check = osd_msg_code; 

    // =============================================================
    // 4. ȭ�� ��� (RGB OSD + HDMI)
    // =============================================================
    
    wire [7:0] vga_r, vga_g, vga_b;

    // (1) RGB ��� (VHDL) �ν��Ͻ�
    // *����: RGB.vhd ������ ������Ʈ �ҽ��� ���ԵǾ� �־�� ��
    RGB u_osd_inst (
        .Din(osd_din),
        .Nblank(cam_href),     // Active Video ��ȣ
        .CLK(clk_pix),         // 25MHz �ȼ� Ŭ��
        .Hsync(cam_href),      // (Ÿ�ֿ̹� �°� HSYNC ����)
        .Vsync(cam_vsync),
        
        // ������ ����
        .msg_code(osd_msg_code),
        .sw(sw),               // SW0, SW2 ��� ���
        .score_c(score_c),
        .score_t(score_t),
        .score_s(score_s),
        
        .R(vga_r),
        .G(vga_g),
        .B(vga_b),
        
        // ��� �� ��
        .x_center(10'd0), .y_center(10'd0), .target_x(10'd0), .target_y(10'd0)
    );

    // (2) HDMI ��ȯ��
    VGA2HDMI u_hdmi_tx (
        .pixclk(clk_pix),
        .clk_TMDS(clk_tmds),
        .VSYNC(cam_vsync),
        .HSYNC(cam_href),     // (���� VGA Ÿ�ֿ̹� �´��� Ȯ�� �ʿ�)
        .ACTIVE(cam_href),
        .red(vga_r),
        .green(vga_g),
        .blue(vga_b),
        .TMDSp(tmds_data_p), .TMDSn(tmds_data_n),
        .TMDSp_clock(tmds_clk_p), .TMDSn_clock(tmds_clk_n)
    );

endmodule